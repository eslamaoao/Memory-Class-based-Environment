package pack;

`include "Transaction.sv"
`include "Sequencer.sv"
`include "Driver.sv"
`include "Monitor.sv"
`include "Scoreboard.sv"
`include "Subscriber.sv"
`include "Env.sv"


endpackage


